
module qsys_led (
	clk_clk,
	led_export,
	sin_export);	

	input		clk_clk;
	output	[15:0]	led_export;
	input	[15:0]	sin_export;
endmodule
